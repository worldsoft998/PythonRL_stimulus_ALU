// sv/uvm_pkg.sv
`ifndef UVM_PKG_SV
`define UVM_PKG_SV
`include "uvm.sv"
`endif
